/*******************************************************************/
/*   ModuleName: tb_PE1  */
/*   Author: Li tianhao    */
/*   Date: 2022/11/1   */
/*   Version: v1.0      */
/********************************************************************/

`timescale 1ns/1ps

module tb_PE1 ();
    
    reg clk;
    reg rstn;
    reg [203:0]  total_blk_i; 
    reg [155:0]  srh_blk_i;
    reg [59:0]  ref_blk_i;
    wire [11:0]  srh_bit_o;
    wire [203:0]  total_blk_o;
    wire [155:0]  srh_blk_o;
    wire [59:0] ref_blk_o;
    wire [7:0] weight_o;

    
    always #10 clk = ~clk;
    
    initial begin
        clk  = 0;
        rstn = 0;
        repeat(10)@(posedge clk);
        rstn = 1;
        repeat(10)@(posedge clk);
        #19
        //case1
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd0};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd0,12'd1,12'd2,12'd3,12'd4};
        #21;
        //case2
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd10};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd0,12'd1,12'd2,12'd3,12'd4};
        #20;
        //case3
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd20};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd0,12'd1,12'd2,12'd3,12'd4};
        #20
        //case4
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd30};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd0,12'd1,12'd2,12'd3,12'd4};
        #20;
        //case5
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd40};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd0,12'd1,12'd2,12'd3,12'd4};
        #20;
        //case6
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd50};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd40,12'd30,12'd20,12'd10,12'd0};
        #20;
        //case7
        srh_blk_i = {12'd1200,12'd1100,12'd1000,12'd900,12'd800,12'd700,12'd600,12'd500,12'd400,12'd300,12'd200,12'd100,12'd60};
        total_blk_i = {12'd180,12'd170,12'd160,12'd150,12'd140,12'd130,12'd120,12'd110,12'd100,12'd90,12'd80,12'd70,12'd60,12'd50,12'd40,12'd30,12'd20,12'd10};
        ref_blk_i = {12'd40,12'd30,12'd20,12'd10,12'd0};
    end
    
    initial begin
        $dumpfile("./build/wave.vcd");  // 指定VCD文件的名字为wave.vcd，仿真信息将记录到此文件
        $dumpvars(0, tb_PE1);  // 指定层次数为0，则tb_code 模块及其下面各层次的�?有信号将被记�?
        #10000$finish;
    end
    
    PE1 u_PE1(
    .clk  (clk),
    .rst_n (rstn),
    .total_blk_i(total_blk_i),
    .srh_blk_i(srh_blk_i),
    .ref_blk_i(ref_blk_i),
    .ref_blk_o(ref_blk_o),
    .srh_bit_o(srh_bit_o),
    .srh_blk_o(srh_blk_o),
    .total_blk_o(total_blk_o),
    .weight_o(weight_o)
    );
    
    
endmodule //tb_PE1
